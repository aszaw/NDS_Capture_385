`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: ECE-Illinois
// Engineer: Zuofu Cheng
// 
// Create Date: 06/08/2023 12:21:05 PM
// Design Name: 
// Module Name: hdmi_text_controller_v1_0_AXI
// Project Name: ECE 385 - hdmi_text_controller
// Target Devices: 
// Tool Versions: 
// Description: 
// This is a modified version of the Vivado template for an AXI4-Lite peripheral,
// rewritten into SystemVerilog for use with ECE 385.
// 
// Dependencies: 
// 
// Revision:
// Revision 0.02 - File modified to be more consistent with generated template
// Revision 11/18 - Made comments less confusing
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


`timescale 1 ns / 1 ps

module hdmi_text_controller_v1_0_AXI #
(

    // Parameters of Axi Slave Bus Interface S_AXI
    // Modify parameters as necessary for access of full VRAM range

    // Width of S_AXI data bus
    parameter integer C_S_AXI_DATA_WIDTH	= 32,
    // Width of S_AXI address bus
    parameter integer C_S_AXI_ADDR_WIDTH	= 16
)
(
    // Users to add ports here
    input logic [9:0] drawX,
    input logic [9:0] drawY,
    output logic inv,
    output logic [10:0] font_addr,
    output logic [11:0] color0,
    output logic [11:0] color1,
    
    // User ports ends

    // Global Clock Signal
    input logic  S_AXI_ACLK,
    // Global Reset Signal. This Signal is Active LOW
    input logic  S_AXI_ARESETN,
    // Write address (issued by master, acceped by Slave)
    input logic [C_S_AXI_ADDR_WIDTH-1 : 0] S_AXI_AWADDR,
    // Write channel Protection type. This signal indicates the
        // privilege and security level of the transaction, and whether
        // the transaction is a data access or an instruction access.
    input logic [2 : 0] S_AXI_AWPROT,
    // Write address valid. This signal indicates that the master signaling
        // valid write address and control information.
    input logic  S_AXI_AWVALID,
    // Write address ready. This signal indicates that the slave is ready
        // to accept an address and associated control signals.
    output logic  S_AXI_AWREADY,
    // Write data (issued by master, acceped by Slave) 
    input logic [C_S_AXI_DATA_WIDTH-1 : 0] S_AXI_WDATA,
    // Write strobes. This signal indicates which byte lanes hold
        // valid data. There is one write strobe bit for each eight
        // bits of the write data bus.    
    input logic [(C_S_AXI_DATA_WIDTH/8)-1 : 0] S_AXI_WSTRB,
    // Write valid. This signal indicates that valid write
        // data and strobes are available.
    input logic  S_AXI_WVALID,
    // Write ready. This signal indicates that the slave
        // can accept the write data.
    output logic  S_AXI_WREADY,
    // Write response. This signal indicates the status
        // of the write transaction.
    output logic [1 : 0] S_AXI_BRESP,
    // Write response valid. This signal indicates that the channel
        // is signaling a valid write response.
    output logic  S_AXI_BVALID,
    // Response ready. This signal indicates that the master
        // can accept a write response.
    input logic  S_AXI_BREADY,
    // Read address (issued by master, acceped by Slave)
    input logic [C_S_AXI_ADDR_WIDTH-1 : 0] S_AXI_ARADDR,
    // Protection type. This signal indicates the privilege
        // and security level of the transaction, and whether the
        // transaction is a data access or an instruction access.
    input logic [2 : 0] S_AXI_ARPROT,
    // Read address valid. This signal indicates that the channel
        // is signaling valid read address and control information.
    input logic  S_AXI_ARVALID,
    // Read address ready. This signal indicates that the slave is
        // ready to accept an address and associated control signals.
    output logic  S_AXI_ARREADY,
    // Read data (issued by slave)
    output logic [C_S_AXI_DATA_WIDTH-1 : 0] S_AXI_RDATA,
    // Read response. This signal indicates the status of the
        // read transfer.
    output logic [1 : 0] S_AXI_RRESP,
    // Read valid. This signal indicates that the channel is
        // signaling the required read data.
    output logic  S_AXI_RVALID,
    // Read ready. This signal indicates that the master can
        // accept the read data and response information.
    input logic  S_AXI_RREADY
);

// AXI4LITE signals
logic  [C_S_AXI_ADDR_WIDTH-1 : 0] 	axi_awaddr;
logic  axi_awready;
logic  axi_wready;
logic  [1 : 0] 	axi_bresp;
logic  axi_bvalid;
logic  [C_S_AXI_ADDR_WIDTH-1 : 0] 	axi_araddr;
logic  axi_arready;
logic  [C_S_AXI_DATA_WIDTH-1 : 0] 	axi_rdata;
logic  [C_S_AXI_DATA_WIDTH-1 : 0] 	axi_wdata;
logic  [1 : 0] 	axi_rresp;
logic  	axi_rvalid;

// Example-specific design signals
// local parameter for addressing 32 bit / 64 bit C_S_AXI_DATA_WIDTH
// ADDR_LSB is used for addressing 32/64 bit registers/memories
// ADDR_LSB = 2 for 32 bits (n downto 2)
// ADDR_LSB = 3 for 64 bits (n downto 3)
localparam integer ADDR_LSB = (C_S_AXI_DATA_WIDTH/32) + 1;
localparam integer OPT_MEM_ADDR_BITS = 9;
//----------------------------------------------
//-- Signals for user logic register space example
//------------------------------------------------
//-- Number of Slave Registers 4
//logic [C_S_AXI_DATA_WIDTH-1:0]	slv_reg0;
//logic [C_S_AXI_DATA_WIDTH-1:0]	slv_reg1;
//logic [C_S_AXI_DATA_WIDTH-1:0]	slv_reg2;
//logic [C_S_AXI_DATA_WIDTH-1:0]	slv_reg3;
//
//Note: the provided Verilog template had the registered declared as above, but in order to give 
//students a hint we have replaced the 4 individual registers with an unpacked array of packed logic. 
//Note that you as the student will still need to extend this to the full register set needed for the lab.
logic [C_S_AXI_DATA_WIDTH-1:0] slv_regs[8];
logic	 slv_reg_rden;
logic	 slv_reg_wren;
logic [C_S_AXI_DATA_WIDTH-1:0]	 reg_data_out;
integer	 byte_index;
logic	 aw_en;

//7.2
logic ReadvramOrPalette; //this is grabing the 14th bit in [13:0] , which is the bit that determines 0 or 2, vram(0) or pallete
logic WriteVramOrPalette;
logic [C_S_AXI_ADDR_WIDTH-1:0] holdval; //holdval is the index of which register it is
logic whichpartofreg;// the last bit of the index, which is 1 or 0, selects which part of the register we want

//assign WriteVramOrPalette = S_AXI_AWADDR[11];   
//assign ReadVramOrPalette = S_AXI_ARADDR[11];
assign WriteVramOrPalette = (S_AXI_AWADDR >= 32'h2000 && S_AXI_AWADDR <= 32'h201F);
assign ReadVramOrPalette = (S_AXI_ARADDR >= 32'h2000 && S_AXI_ARADDR <= 32'h201F);


// I/O Connections assignments

assign S_AXI_AWREADY = axi_awready;
assign S_AXI_WREADY	= axi_wready;
assign S_AXI_BRESP	= axi_bresp;
assign S_AXI_BVALID	= axi_bvalid;
assign S_AXI_ARREADY = axi_arready;
//assign S_AXI_WDATA = axi_wdata;
assign S_AXI_RDATA = axi_rdata;
assign S_AXI_RRESP	= axi_rresp;
assign S_AXI_RVALID	= axi_rvalid;

// Implement axi_awready generation
// axi_awready is asserted for one S_AXI_ACLK clock cycle when both
// S_AXI_AWVALID and S_AXI_WVALID are asserted. axi_awready is
// de-asserted when reset is low.

always_ff @( posedge S_AXI_ACLK )
begin
  if ( S_AXI_ARESETN == 1'b0 )
    begin
      axi_awready <= 1'b0;
      aw_en <= 1'b1;
    end 
  else
    begin    
      if (~axi_awready && S_AXI_AWVALID && S_AXI_WVALID && aw_en)
        begin
          // slave is ready to accept write address when 
          // there is a valid write address and write data
          // on the write address and data bus. This design 
          // expects no outstanding transactions. 
          axi_awready <= 1'b1;
          aw_en <= 1'b0;
        end
        else if (S_AXI_BREADY && axi_bvalid)
            begin
              aw_en <= 1'b1;
              axi_awready <= 1'b0;
            end
      else           
        begin
          axi_awready <= 1'b0;
        end
    end 
end       

// Implement axi_awaddr latching
// This process is used to latch the address when both 
// S_AXI_AWVALID and S_AXI_WVALID are valid. 

always_ff @( posedge S_AXI_ACLK )
begin
  if ( S_AXI_ARESETN == 1'b0 )
    begin
      axi_awaddr <= 0;
    end 
  else
    begin    
      if (~axi_awready && S_AXI_AWVALID && S_AXI_WVALID && aw_en)
        begin
          // Write Address latching 
          axi_awaddr <= S_AXI_AWADDR;
        end
    end 
end       

// Implement axi_wready generation
// axi_wready is asserted for one S_AXI_ACLK clock cycle when both
// S_AXI_AWVALID and S_AXI_WVALID are asserted. axi_wready is 
// de-asserted when reset is low. 

always_ff @( posedge S_AXI_ACLK )
begin
  if ( S_AXI_ARESETN == 1'b0 )
    begin
      axi_wready <= 1'b0;
    end 
  else
    begin    
      if (~axi_wready && S_AXI_WVALID && S_AXI_AWVALID && aw_en )
        begin
          // slave is ready to accept write data when 
          // there is a valid write address and write data
          // on the write address and data bus. This design 
          // expects no outstanding transactions. 
          axi_wready <= 1'b1;
        end
      else
        begin
          axi_wready <= 1'b0;
        end
    end 
end       

// Implement memory mapped register select and write logic generation
// The write data is accepted and written to memory mapped registers when
// axi_awready, S_AXI_WVALID, axi_wready and S_AXI_WVALID are asserted. Write strobes are used to
// select byte enables of slave registers while writing.
// These registers are cleared when reset (active low) is applied.
// Slave register write enable is asserted when valid address and data are available
// and the slave is ready to accept the write address and write data.
 
assign slv_reg_wren = axi_wready && S_AXI_WVALID && axi_awready && S_AXI_AWVALID;
assign slv_reg_rden = axi_arready && S_AXI_ARVALID && ~axi_rvalid;

// 7.2
logic [3:0] strobe;
logic [15:0] findaddr;
logic [31:0] dataAin;


always_ff @( posedge S_AXI_ACLK )
    begin
//         if ( S_AXI_ARESETN == 1'b0 )
//            begin
//                 axi_rdata <= 16'h0000;
//                 for (integer i = 0; i < 9; i++) begin
//                    slv_regs[i] <= 0;
//                 end
//            end
            //vram write
              if(slv_reg_wren == 1 && WriteVramOrPalette == 1'b0)begin 
                findaddr <= S_AXI_AWADDR[ADDR_LSB+OPT_MEM_ADDR_BITS:ADDR_LSB]; 
                strobe <= S_AXI_WSTRB;
                dataAin <= S_AXI_WDATA;
               end
              //vram read
               else if (slv_reg_rden && ReadVramOrPalette == 1'b0)begin
                       findaddr <= axi_araddr[ADDR_LSB+OPT_MEM_ADDR_BITS:ADDR_LSB];
                       strobe <= 4'b0000;
                       axi_rdata <= dataAout;
               end
               //palette reg B write
               else if( slv_reg_wren == 1 && WriteVramOrPalette == 1'b1 )begin 
                    for (byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1) begin
                        if (S_AXI_WSTRB[byte_index]) begin
                            slv_regs[axi_awaddr[4:2]][(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +:8];
                        end else begin
                             slv_regs[axi_awaddr[4:2]][(byte_index*8) +: 8] <= slv_regs[axi_awaddr[4:2]][(byte_index*8) +: 8];
                        end
                    end
               end 
               //pallete reg B read
               else if (slv_reg_rden == 1 && ReadVramOrPalette == 1'b1 )begin
                    axi_rdata <= slv_regs[axi_araddr[4:2]];
               end
    end    


// Implement write response logic generation
// The write response and response valid signals are asserted by the slave 
// when axi_wready, S_AXI_WVALID, axi_wready and S_AXI_WVALID are asserted.  
// This marks the acceptance of address and indicates the status of 
// write transaction.

always_ff @( posedge S_AXI_ACLK )
begin
  if ( S_AXI_ARESETN == 1'b0 )
    begin
      axi_bvalid  <= 1'b0;
      axi_bresp   <= 2'b0;
    end 
  else
    begin    
      if (axi_awready && S_AXI_AWVALID && ~axi_bvalid && axi_wready && S_AXI_WVALID)
        begin
          // indicates a valid write response is available
          axi_bvalid <= 1'b1;
          axi_bresp  <= 2'b0; // 'OKAY' response 
        end                   // work error responses in future
      else
        begin
          if (S_AXI_BREADY && axi_bvalid) 
            //check if bready is asserted while bvalid is high) 
            //(there is a possibility that bready is always asserted high)   
            begin
              axi_bvalid <= 1'b0; 
            end  
        end
    end
end   

// Implement axi_arready generation
// axi_arready is asserted for one S_AXI_ACLK clock cycle when
// S_AXI_ARVALID is asserted. axi_awready is 
// de-asserted when reset (active low) is asserted. 
// The read address is also latched when S_AXI_ARVALID is 
// asserted. axi_araddr is reset to zero on reset assertion.

always_ff @( posedge S_AXI_ACLK )
begin
  if ( S_AXI_ARESETN == 1'b0 )
    begin
      axi_arready <= 1'b0;
      axi_araddr  <= 32'b0;
    end 
  else
    begin    
      if (~axi_arready && S_AXI_ARVALID)
        begin
          // indicates that the slave has acceped the valid read address
          axi_arready <= 1'b1;
          // Read address latching
          axi_araddr  <= S_AXI_ARADDR;
        end
      else
        begin
          axi_arready <= 1'b0;
        end
    end 
end       

// Implement axi_arvalid generation
// axi_rvalid is asserted for one S_AXI_ACLK clock cycle when both 
// S_AXI_ARVALID and axi_arready are asserted. The slave registers 
// data are available on the axi_rdata bus at this instance. The 
// assertion of axi_rvalid marks the validity of read data on the 
// bus and axi_rresp indicates the status of read transaction.axi_rvalid 
// is deasserted on reset (active low). axi_rresp and axi_rdata are 
// cleared to zero on reset (active low).  
always_ff @( posedge S_AXI_ACLK )
begin
  if ( S_AXI_ARESETN == 1'b0 )
    begin
      axi_rdata <= 0;
      axi_rvalid <= 0;
      axi_rresp  <= 0;
    end 
  else
    begin    
      if (axi_arready && S_AXI_ARVALID && ~axi_rvalid)
        begin
          // Valid read data is available at the read data bus
          axi_rvalid <= 1'b1;
          axi_rresp  <= 2'b0; // 'OKAY' response
        end   
      else if (axi_rvalid && S_AXI_RREADY)
        begin
          // Read data is accepted by the master
          axi_rvalid <= 1'b0;
        end                
    end
end    

// Implement memory mapped register select and read logic generation
// Slave register read enable is asserted when valid address is available
// and the slave is ready to accept the read address.

//assign slv_reg_rden = axi_arready & S_AXI_ARVALID & ~axi_rvalid;

//always_comb
//begin
//      // Address decoding for reading registers
//     reg_data_out = slv_regs[axi_araddr[ADDR_LSB+OPT_MEM_ADDR_BITS:ADDR_LSB]];
//end

// Output register or memory read data
//always_ff @( posedge S_AXI_ACLK )
//begin
//  if ( S_AXI_ARESETN == 1'b0 )
//    begin
//      axi_rdata  <= 0;
//    end 
//  else
//    begin    
//      // When there is a valid read address (S_AXI_ARVALID) with 
//      // acceptance of read address by the slave (axi_arready), 
//      // output the read dada 
//      if (slv_reg_rden)
//        begin
//          axi_rdata <= reg_data_out;     // register read data
//        end   
//    end
//end    

logic [31:0] dummy;
logic [31:0] dataAout;
logic [15:0] addrb;
logic [15:0] hold;

//assign holdval = drawX[9:3] + (drawY[9:4]*80);
logic [9:0] col, row;
assign col = drawX >> 3;
assign row = drawY >> 4;
//assign hold = row * 80 + (col);
assign hold =  drawX[9:3] + (drawY[9:4]*80);
assign whichpartofreg = hold[0];
assign addrb = hold >> 1;

logic [31:0]outputReg;

//assign addrb = holdval >> 1;

blk_mem_gen_0 ram(.addra(findaddr), //findaddr
                .clka(S_AXI_ACLK), 
                .dina(dataAin), 
                .douta(dataAout), 
                .ena(1'b1), 
                .wea(strobe), //S_AXI_WDATA//S_AXI_RDATA
                
                .addrb(addrb), 
                .clkb(S_AXI_ACLK), 
                .dinb(dummy), 
                .doutb(outputReg), 
                .enb(1'b1), 
                .web(4'h0000));
                
// Add user logic here

logic [7:0] char_code;
logic [3:0] fg_idx;
logic [3:0] bg_idx;

always_comb begin
        //WhaStIsInTheReg <= slv_regs[(DrawY/16)*20+ DrawX/32];//This line grabs the data inside of the specific register
        //WhatPartOfReg <= WhatIsInTheReg[((DrawX % 32)/8)*8 +: 8];//What part(which 8 bits do we want)
        
        if(whichpartofreg == 1'b1)begin
            char_code = outputReg[31:24];
            fg_idx = outputReg[23:20];
            bg_idx = outputReg[19:16];
        end
        else begin
            char_code = outputReg[15:8];
            fg_idx = outputReg[7:4];
            bg_idx = outputReg[3:0];
        end
        
        inv = char_code[7];
        font_addr = (char_code[6:0] * 16) + (drawY[3:0]); // output this to fontrom to get the data
        if(fg_idx[0] == 1'b1)begin
            color1 = slv_regs[fg_idx >> 1][24:13];
        end
        else begin
            color1 =  slv_regs[fg_idx >> 1][12:1];
        end
        
        if(bg_idx[0] == 1'b1)begin
            color0 =  slv_regs[bg_idx >> 1][24:13];
        end
        else begin
            color0 =  slv_regs[bg_idx >> 1][12:1];
        end
        
end


//logic [9:0] row, col;
//logic [11:0] regis;
//logic [1:0] char;
//logic [7:0] char_code;

//always_comb
//begin 
//    row  = drawY >> 4;
//    col = drawX >> 2;
    
//    regis = row * 20 + (col >>2 );
//    char = col[1:0];
//    outputReg = slv_regs[600];
//    case(char)
//        2'b00: char_code = slv_regs[regis][7:0];
//        2'b01: char_code = slv_regs[regis][15:8];
//        2'b10: char_code = slv_regs[regis][23:16];
//        2'b11: char_code = slv_regs[regis][31:24];
//    endcase
//   // inv = char_code[7];
//    font_addr = (char_code[6:0] << 4) + drawY[3:0];
//end

// User logic ends

endmodule